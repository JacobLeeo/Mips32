module EX(
  input  [7:0]  io_inFromD_iSK,
  input  [2:0]  io_inFromD_iK,
  input  [31:0] io_inFromD_source1,
  input  [31:0] io_inFromD_source2,
  input  [4:0]  io_inFromD_rWAddr,
  input         io_inFromD_rWEn,
  output [4:0]  io_outToD_rWAddrO,
  output        io_outToD_rWEnO,
  output [31:0] io_outToD_rWDataO
);
  wire [31:0] _logicResult_T = io_inFromD_source1 | io_inFromD_source2; // @[EX.scala 30:47]
  wire [31:0] logicResult = 8'h25 == io_inFromD_iSK ? _logicResult_T : 32'h0; // @[EX.scala 28:28 30:25]
  assign io_outToD_rWAddrO = io_inFromD_rWAddr; // @[EX.scala 21:23]
  assign io_outToD_rWEnO = io_inFromD_rWEn; // @[EX.scala 22:21]
  assign io_outToD_rWDataO = 3'h1 == io_inFromD_iK ? logicResult : 32'h0; // @[EX.scala 24:23 35:27 37:31]
endmodule
module DbtEXMEM(
  input         clock,
  input  [4:0]  io_inFromEX_rWAddrO,
  input         io_inFromEX_rWEnO,
  input  [31:0] io_inFromEX_rWDataO,
  output [4:0]  io_outToMEM_rWAddrO,
  output        io_outToMEM_rWEnO,
  output [31:0] io_outToMEM_rWDataO
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] rWAddr; // @[DbtEXMEM.scala 19:25]
  reg  rWEn; // @[DbtEXMEM.scala 20:23]
  reg [31:0] rWData; // @[DbtEXMEM.scala 21:25]
  assign io_outToMEM_rWAddrO = rWAddr; // @[DbtEXMEM.scala 23:25]
  assign io_outToMEM_rWEnO = rWEn; // @[DbtEXMEM.scala 24:23]
  assign io_outToMEM_rWDataO = rWData; // @[DbtEXMEM.scala 25:25]
  always @(posedge clock) begin
    rWAddr <= io_inFromEX_rWAddrO; // @[DbtEXMEM.scala 19:25]
    rWEn <= io_inFromEX_rWEnO; // @[DbtEXMEM.scala 20:23]
    rWData <= io_inFromEX_rWDataO; // @[DbtEXMEM.scala 21:25]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rWAddr = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  rWEn = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  rWData = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EXTop(
  input         clock,
  input         reset,
  input  [7:0]  io_inFromID_iSK,
  input  [2:0]  io_inFromID_iK,
  input  [31:0] io_inFromID_source1,
  input  [31:0] io_inFromID_source2,
  input  [4:0]  io_inFromID_rWAddr,
  input         io_inFromID_rWEn,
  output [4:0]  io_outToMEM_rWAddrO,
  output        io_outToMEM_rWEnO,
  output [31:0] io_outToMEM_rWDataO
);
  wire [7:0] ex_io_inFromD_iSK; // @[EXTop.scala 13:20]
  wire [2:0] ex_io_inFromD_iK; // @[EXTop.scala 13:20]
  wire [31:0] ex_io_inFromD_source1; // @[EXTop.scala 13:20]
  wire [31:0] ex_io_inFromD_source2; // @[EXTop.scala 13:20]
  wire [4:0] ex_io_inFromD_rWAddr; // @[EXTop.scala 13:20]
  wire  ex_io_inFromD_rWEn; // @[EXTop.scala 13:20]
  wire [4:0] ex_io_outToD_rWAddrO; // @[EXTop.scala 13:20]
  wire  ex_io_outToD_rWEnO; // @[EXTop.scala 13:20]
  wire [31:0] ex_io_outToD_rWDataO; // @[EXTop.scala 13:20]
  wire  d_clock; // @[EXTop.scala 14:19]
  wire [4:0] d_io_inFromEX_rWAddrO; // @[EXTop.scala 14:19]
  wire  d_io_inFromEX_rWEnO; // @[EXTop.scala 14:19]
  wire [31:0] d_io_inFromEX_rWDataO; // @[EXTop.scala 14:19]
  wire [4:0] d_io_outToMEM_rWAddrO; // @[EXTop.scala 14:19]
  wire  d_io_outToMEM_rWEnO; // @[EXTop.scala 14:19]
  wire [31:0] d_io_outToMEM_rWDataO; // @[EXTop.scala 14:19]
  EX ex ( // @[EXTop.scala 13:20]
    .io_inFromD_iSK(ex_io_inFromD_iSK),
    .io_inFromD_iK(ex_io_inFromD_iK),
    .io_inFromD_source1(ex_io_inFromD_source1),
    .io_inFromD_source2(ex_io_inFromD_source2),
    .io_inFromD_rWAddr(ex_io_inFromD_rWAddr),
    .io_inFromD_rWEn(ex_io_inFromD_rWEn),
    .io_outToD_rWAddrO(ex_io_outToD_rWAddrO),
    .io_outToD_rWEnO(ex_io_outToD_rWEnO),
    .io_outToD_rWDataO(ex_io_outToD_rWDataO)
  );
  DbtEXMEM d ( // @[EXTop.scala 14:19]
    .clock(d_clock),
    .io_inFromEX_rWAddrO(d_io_inFromEX_rWAddrO),
    .io_inFromEX_rWEnO(d_io_inFromEX_rWEnO),
    .io_inFromEX_rWDataO(d_io_inFromEX_rWDataO),
    .io_outToMEM_rWAddrO(d_io_outToMEM_rWAddrO),
    .io_outToMEM_rWEnO(d_io_outToMEM_rWEnO),
    .io_outToMEM_rWDataO(d_io_outToMEM_rWDataO)
  );
  assign io_outToMEM_rWAddrO = d_io_outToMEM_rWAddrO; // @[EXTop.scala 18:19]
  assign io_outToMEM_rWEnO = d_io_outToMEM_rWEnO; // @[EXTop.scala 18:19]
  assign io_outToMEM_rWDataO = d_io_outToMEM_rWDataO; // @[EXTop.scala 18:19]
  assign ex_io_inFromD_iSK = io_inFromID_iSK; // @[EXTop.scala 16:19]
  assign ex_io_inFromD_iK = io_inFromID_iK; // @[EXTop.scala 16:19]
  assign ex_io_inFromD_source1 = io_inFromID_source1; // @[EXTop.scala 16:19]
  assign ex_io_inFromD_source2 = io_inFromID_source2; // @[EXTop.scala 16:19]
  assign ex_io_inFromD_rWAddr = io_inFromID_rWAddr; // @[EXTop.scala 16:19]
  assign ex_io_inFromD_rWEn = io_inFromID_rWEn; // @[EXTop.scala 16:19]
  assign d_clock = clock;
  assign d_io_inFromEX_rWAddrO = ex_io_outToD_rWAddrO; // @[EXTop.scala 17:18]
  assign d_io_inFromEX_rWEnO = ex_io_outToD_rWEnO; // @[EXTop.scala 17:18]
  assign d_io_inFromEX_rWDataO = ex_io_outToD_rWDataO; // @[EXTop.scala 17:18]
endmodule
